package fifo_tb_pkg;

    `include "transaction_base.sv"
    `include "component.sv"
    `include "fifo_transaction.sv"
    `include "fifo_generator.sv"
    `include "fifo_driver.sv"
    `include "fifo_monitor.sv"
    `include "environment.sv"  
    
endpackage
  